-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition
-- Created on Sun Jul 27 15:12:23 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachineEditor IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        din : IN STD_LOGIC := '0';
        den : IN STD_LOGIC := '0';
        dvalid : IN STD_LOGIC := '0';
        dmatch : IN STD_LOGIC := '0';
        sync : OUT STD_LOGIC
    );
END StateMachineEditor;

ARCHITECTURE BEHAVIOR OF StateMachineEditor IS
    TYPE type_fstate IS (NOT_MATCHING,MATCHING,MATCHING_END,SYNC);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,din,den,dvalid,dmatch)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= NOT_MATCHING;
            sync <= '0';
        ELSE
            sync <= '0';
            CASE fstate IS
                WHEN NOT_MATCHING =>
                    IF ((((den = '1') AND (din = dmatch)) AND (dvalid = '1'))) THEN
                        reg_fstate <= MATCHING;
                    ELSE
                        reg_fstate <= NOT_MATCHING;
                    END IF;

                    sync <= '0';
                WHEN MATCHING =>
                    IF (((den = '1') AND ((din /= dmatch) OR (dvalid = '0')))) THEN
                        reg_fstate <= MATCHING_END;
                    ELSE
                        reg_fstate <= MATCHING;
                    END IF;

                    sync <= '0';
                WHEN MATCHING_END =>
                    IF ((((den = '1') AND (din /= dmatch)) AND (dvalid = '1'))) THEN
                        reg_fstate <= SYNC;
                    ELSIF (((den = '0') OR ((dmatch = din) AND (dvalid = '1')))) THEN
                        reg_fstate <= MATCHING_END;
                    ELSE
                        reg_fstate <= NOT_MATCHING;
                    END IF;

                    sync <= '0';
                WHEN SYNC =>
                    reg_fstate <= NOT_MATCHING;

                    sync <= '1';
                WHEN OTHERS => 
                    sync <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
